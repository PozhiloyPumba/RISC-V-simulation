module V
(
	input clk,
	input rst
);

RV32 RV32(.clk(clk), .rst(rst));

endmodule