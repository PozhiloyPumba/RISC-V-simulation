module CU
(
    
);
    
endmodule