module DECODER
(
    
);
    
endmodule