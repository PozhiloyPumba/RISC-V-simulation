module ALU
(
    
);


endmodule